module E#(


    
)