module hazard(
    //FORWARDING   
    input Rs1E
    input Rs2E

)

endmodule