module Hazard(
    //FORWARDING   
    input Rs1E
    input Rs2E

)

endmodule